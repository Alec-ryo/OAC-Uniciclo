library ieee; 
use ieee.std_logic_1164.all; 

package xregs_pkg is

type registradores is array (31 downto 0) of std_logic_vector(31 downto 0);

end xregs_pkg;