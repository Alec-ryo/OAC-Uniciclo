package imm_pkg is 

type FORMAT_RV is ( R_type, I_type, S_type, SB_type, UJ_type, U_type );

end imm_pkg;
