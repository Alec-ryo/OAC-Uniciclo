package rv_pkg is 

type ULA_OP is ( ADD_OP, SUB_OP, AND_OP, OR_OP, NOR_OP,
					  XOR_OP, SLL_OP, SRL_OP, SRA_OP, SLT_OP,
					  SLTU_OP, SGE_OP, SGEU_OP, SEQ_OP, SNE_OP
);

end rv_pkg;
